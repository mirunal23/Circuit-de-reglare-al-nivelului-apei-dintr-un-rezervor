** Profile: "SCHEMATIC1-montecarlo_timp"  [ C:\Miruna\PROIECT_ORCAD\Proiect-PSpiceFiles\SCHEMATIC1\montecarlo_timp.sim ] 

** Creating circuit file "montecarlo_timp.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../dportocala.lib" 
* From [PSPICE NETLIST] section of C:\SPB_Data\cdssetup\OrCAD_PSpice\22.1.0\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 10ms 0 
.MC 50 TRAN V([OUT]) YMAX OUTPUT ALL SEED=200 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
