** Profile: "SCHEMATIC1-Worst_Case"  [ C:\Miruna\PROIECT_ORCAD\proiect-pspicefiles\schematic1\worst_case.sim ] 

** Creating circuit file "Worst_Case.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../dportocala.lib" 
* From [PSPICE NETLIST] section of C:\SPB_Data\cdssetup\OrCAD_PSpice\22.1.0\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.DC LIN PARAM r 35k 15k 100 
.WCASE DC V([OUT]) YMAX VARY BOTH  HI 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
