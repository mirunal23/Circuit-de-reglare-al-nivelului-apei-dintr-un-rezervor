** Profile: "SCHEMATIC1-dioda"  [ C:\Miruna\PROIECT_ORCAD\Proiect-PSpiceFiles\SCHEMATIC1\dioda.sim ] 

** Creating circuit file "dioda.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../dportocala.lib" 
* From [PSPICE NETLIST] section of C:\SPB_Data\cdssetup\OrCAD_PSpice\22.1.0\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.DC LIN V_V3 0 3 0.1 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
